// This file contains a pareto-optimal circuit with respect to power and the fault-resilince parameter p_fault which is defined as:
// "For all input vectors, the ratio of the no. of faults observable at the POs to the no. of total possible faults in the circuit".
// This code is part of the ReCkt library (https://github.com/umar-afzaal/ReCkt) distributed under The MIT License.
// When used, please cite the following article(s):
// U. Afzaal, A.S. Hassan, M. Usman and J.A. Lee, "On the Evolutionary Synthesis of Increased Fault-resilience Arithmetic Circuits".

// p_fault = 77.1 %    (Lower is better)
// gates = 26.0
// levels = 9
// area = 36.32    (For MCNC library relative to nand2)
// power = 102.0 uW    (Berkely-SIS for MCNC library @ Vdd=5V and 20 MHz clock)
// delay = 14.8 ns    (Berkely-ABC for MCNC library)
// PDP = 1.5096e-12 J

// Pin mapping:
// {n0, n1, n2, n3} = A[3:0]
// {n4, n5, n6, n7} = B[3:0]
// {n25, n23, n20, n18, n34} = O[4:0]

module addr4u_power_11 (
n0, n1, n2, n3, n4, n5, n6, n7, 
n25, n23, n20, n18, n34
);

input n0, n1, n2, n3, n4, n5, n6, n7;
output n25, n23, n20, n18, n34;
wire n29, n13, n30, n24, n9, n14, n16, n8, n22, n15, n10, n31, n26, n19, n21, n33, n27, n11, n28, n12, 
n17;

xor (n8, n4, n0);
nand (n9, n4, n0);
nand (n10, n5, n1);
nand (n11, n6, n2);
nor (n12, n7, n3);
xor (n13, n6, n2);
and (n14, n7, n3);
xor (n15, n5, n1);
nor (n16, n12, n14);
nand (n17, n13, n14);
xor (n18, n13, n14);
nand (n19, n17, n11);
xor (n20, n15, n19);
nand (n21, n15, n19);
nand (n22, n21, n10);
xor (n23, n8, n22);
nand (n24, n8, n22);
nand (n25, n24, n9);
xor (n26, n20, n20);
xor (n27, n20, n20);
and (n28, n27, n26);
xor (n29, n26, n27);
nand (n30, n16, n16);
and (n31, n28, n29);
and (n33, n29, n31);
nor (n34, n33, n30);

endmodule